`timescale 1ns/ 1ps

module fc_weights_memory(
    input wire clk,
    input wire rst,
    input wire start,
    input wire [5: 0] input_pixel_addr,
    input wire [4: 0] output_pixel_addr,
    output reg signed [15: 0] w,
    output reg signed [31: 0] b,
    output reg ready
);
    reg signed [15: 0] weights [0: 31][0: 59];
    reg signed [31: 0] biases [0: 31];

    initial begin
        weights[ 0][0]<=-192;  weights[ 0][1]<= 153;  weights[ 0][2]<= 109;  weights[ 0][3]<= -32;  weights[ 0][4]<= 198;  weights[ 0][5]<=  -2;  weights[ 0][6]<=-271;  weights[ 0][7]<= 149;  weights[ 0][8]<=  73;  weights[ 0][9]<= -33;  weights[ 0][10]<=  84;  weights[ 0][11]<= 100;  weights[ 0][12]<=-117;  weights[ 0][13]<=  76;  weights[ 0][14]<=-114;  weights[ 0][15]<=  60;  weights[ 0][16]<=  29;  weights[ 0][17]<=  85;  weights[ 0][18]<= 131;  weights[ 0][19]<= 131;  weights[ 0][20]<= 176;  weights[ 0][21]<= 166;  weights[ 0][22]<= 128;  weights[ 0][23]<=-139;  weights[ 0][24]<= 154;  weights[ 0][25]<=  53;  weights[ 0][26]<=-144;  weights[ 0][27]<=-149;  weights[ 0][28]<= -80;  weights[ 0][29]<=-102;  weights[ 0][30]<=-221;  weights[ 0][31]<=  35;  weights[ 0][32]<= 157;  weights[ 0][33]<=-273;  weights[ 0][34]<= -52;  weights[ 0][35]<=  76;  weights[ 0][36]<= -52;  weights[ 0][37]<=-122;  weights[ 0][38]<= 235;  weights[ 0][39]<=  88;  weights[ 0][40]<=-155;  weights[ 0][41]<=-164;  weights[ 0][42]<= -26;  weights[ 0][43]<=-150;  weights[ 0][44]<=  25;  weights[ 0][45]<=  25;  weights[ 0][46]<=-148;  weights[ 0][47]<=  15;  weights[ 0][48]<=-113;  weights[ 0][49]<=-152;  weights[ 0][50]<= 163;  weights[ 0][51]<=  35;  weights[ 0][52]<=-168;  weights[ 0][53]<= 114;  weights[ 0][54]<= -91;  weights[ 0][55]<=-112;  weights[ 0][56]<=  81;  weights[ 0][57]<= -90;  weights[ 0][58]<=-147;  weights[ 0][59]<=-166;  
        weights[ 1][0]<= 128;  weights[ 1][1]<= 263;  weights[ 1][2]<= -42;  weights[ 1][3]<= 175;  weights[ 1][4]<=-135;  weights[ 1][5]<=-204;  weights[ 1][6]<= -11;  weights[ 1][7]<=  18;  weights[ 1][8]<= 226;  weights[ 1][9]<= -85;  weights[ 1][10]<= 223;  weights[ 1][11]<=  90;  weights[ 1][12]<=-105;  weights[ 1][13]<=  68;  weights[ 1][14]<=  91;  weights[ 1][15]<=-198;  weights[ 1][16]<=-317;  weights[ 1][17]<=  20;  weights[ 1][18]<= 172;  weights[ 1][19]<=-113;  weights[ 1][20]<= 157;  weights[ 1][21]<= -38;  weights[ 1][22]<= -52;  weights[ 1][23]<=-120;  weights[ 1][24]<=-131;  weights[ 1][25]<= 273;  weights[ 1][26]<=-191;  weights[ 1][27]<=-138;  weights[ 1][28]<=  89;  weights[ 1][29]<=  89;  weights[ 1][30]<=-135;  weights[ 1][31]<= 194;  weights[ 1][32]<=-123;  weights[ 1][33]<= -97;  weights[ 1][34]<=  80;  weights[ 1][35]<= 186;  weights[ 1][36]<=  60;  weights[ 1][37]<= 137;  weights[ 1][38]<= -93;  weights[ 1][39]<= -94;  weights[ 1][40]<=  -1;  weights[ 1][41]<=-182;  weights[ 1][42]<=  38;  weights[ 1][43]<= 126;  weights[ 1][44]<=-103;  weights[ 1][45]<=-141;  weights[ 1][46]<= -27;  weights[ 1][47]<= -11;  weights[ 1][48]<= -45;  weights[ 1][49]<=  34;  weights[ 1][50]<= 110;  weights[ 1][51]<=-168;  weights[ 1][52]<= 136;  weights[ 1][53]<= -37;  weights[ 1][54]<=-168;  weights[ 1][55]<= -80;  weights[ 1][56]<= -13;  weights[ 1][57]<= -74;  weights[ 1][58]<=  55;  weights[ 1][59]<=-109;  
        weights[ 2][0]<= -94;  weights[ 2][1]<=-146;  weights[ 2][2]<= 138;  weights[ 2][3]<= 157;  weights[ 2][4]<= -25;  weights[ 2][5]<=-132;  weights[ 2][6]<= 208;  weights[ 2][7]<= -67;  weights[ 2][8]<= -51;  weights[ 2][9]<=-177;  weights[ 2][10]<=  24;  weights[ 2][11]<=  76;  weights[ 2][12]<= 111;  weights[ 2][13]<=-113;  weights[ 2][14]<=  22;  weights[ 2][15]<=  24;  weights[ 2][16]<= 168;  weights[ 2][17]<= 178;  weights[ 2][18]<= 113;  weights[ 2][19]<= -26;  weights[ 2][20]<= 161;  weights[ 2][21]<= 204;  weights[ 2][22]<=   1;  weights[ 2][23]<=-115;  weights[ 2][24]<=  -1;  weights[ 2][25]<= 198;  weights[ 2][26]<=  57;  weights[ 2][27]<=  59;  weights[ 2][28]<=-210;  weights[ 2][29]<= 123;  weights[ 2][30]<= 148;  weights[ 2][31]<= 196;  weights[ 2][32]<=  26;  weights[ 2][33]<=  -2;  weights[ 2][34]<= 166;  weights[ 2][35]<= 122;  weights[ 2][36]<= 106;  weights[ 2][37]<=  94;  weights[ 2][38]<=-223;  weights[ 2][39]<=  -3;  weights[ 2][40]<=-193;  weights[ 2][41]<=  21;  weights[ 2][42]<= 160;  weights[ 2][43]<=-132;  weights[ 2][44]<= -81;  weights[ 2][45]<= 120;  weights[ 2][46]<= 167;  weights[ 2][47]<= 275;  weights[ 2][48]<=-197;  weights[ 2][49]<=-153;  weights[ 2][50]<= -17;  weights[ 2][51]<=-109;  weights[ 2][52]<=  32;  weights[ 2][53]<=-167;  weights[ 2][54]<=  66;  weights[ 2][55]<=-187;  weights[ 2][56]<=  80;  weights[ 2][57]<=  75;  weights[ 2][58]<=-107;  weights[ 2][59]<= -83;  
        weights[ 3][0]<=   9;  weights[ 3][1]<= 203;  weights[ 3][2]<= 135;  weights[ 3][3]<= 143;  weights[ 3][4]<=-210;  weights[ 3][5]<= -61;  weights[ 3][6]<=  51;  weights[ 3][7]<=  35;  weights[ 3][8]<=  84;  weights[ 3][9]<=  40;  weights[ 3][10]<= -55;  weights[ 3][11]<= 114;  weights[ 3][12]<= 123;  weights[ 3][13]<=  25;  weights[ 3][14]<= 205;  weights[ 3][15]<=  36;  weights[ 3][16]<= 202;  weights[ 3][17]<=-123;  weights[ 3][18]<=-226;  weights[ 3][19]<=  19;  weights[ 3][20]<= 110;  weights[ 3][21]<= 158;  weights[ 3][22]<= 228;  weights[ 3][23]<= -85;  weights[ 3][24]<=-171;  weights[ 3][25]<= 152;  weights[ 3][26]<= -64;  weights[ 3][27]<=   1;  weights[ 3][28]<= -29;  weights[ 3][29]<= -29;  weights[ 3][30]<= 145;  weights[ 3][31]<=  70;  weights[ 3][32]<=-181;  weights[ 3][33]<= -55;  weights[ 3][34]<=-238;  weights[ 3][35]<=  24;  weights[ 3][36]<=-215;  weights[ 3][37]<= 169;  weights[ 3][38]<=-254;  weights[ 3][39]<= 126;  weights[ 3][40]<=   5;  weights[ 3][41]<= -12;  weights[ 3][42]<=   1;  weights[ 3][43]<= 222;  weights[ 3][44]<=  40;  weights[ 3][45]<=-120;  weights[ 3][46]<=  55;  weights[ 3][47]<=-120;  weights[ 3][48]<=   3;  weights[ 3][49]<=  66;  weights[ 3][50]<=-212;  weights[ 3][51]<= -72;  weights[ 3][52]<=  80;  weights[ 3][53]<=  47;  weights[ 3][54]<=-145;  weights[ 3][55]<= 133;  weights[ 3][56]<=   3;  weights[ 3][57]<= -67;  weights[ 3][58]<= -37;  weights[ 3][59]<= 165;  
        weights[ 4][0]<=   6;  weights[ 4][1]<= -93;  weights[ 4][2]<=-217;  weights[ 4][3]<=-127;  weights[ 4][4]<=-136;  weights[ 4][5]<=-197;  weights[ 4][6]<= 200;  weights[ 4][7]<= -45;  weights[ 4][8]<=  42;  weights[ 4][9]<=  11;  weights[ 4][10]<=-162;  weights[ 4][11]<= -70;  weights[ 4][12]<= -17;  weights[ 4][13]<= 273;  weights[ 4][14]<=  55;  weights[ 4][15]<=-106;  weights[ 4][16]<= 200;  weights[ 4][17]<=  34;  weights[ 4][18]<= -20;  weights[ 4][19]<=  16;  weights[ 4][20]<= 228;  weights[ 4][21]<= 169;  weights[ 4][22]<=  52;  weights[ 4][23]<= 115;  weights[ 4][24]<= 252;  weights[ 4][25]<= -68;  weights[ 4][26]<= -45;  weights[ 4][27]<=  87;  weights[ 4][28]<=-207;  weights[ 4][29]<=-142;  weights[ 4][30]<=-117;  weights[ 4][31]<= -53;  weights[ 4][32]<=  80;  weights[ 4][33]<= 255;  weights[ 4][34]<= 145;  weights[ 4][35]<= -96;  weights[ 4][36]<=-215;  weights[ 4][37]<= 208;  weights[ 4][38]<=  -5;  weights[ 4][39]<=  56;  weights[ 4][40]<= 187;  weights[ 4][41]<=-225;  weights[ 4][42]<=-105;  weights[ 4][43]<=   0;  weights[ 4][44]<=  80;  weights[ 4][45]<=  -4;  weights[ 4][46]<= 102;  weights[ 4][47]<=-208;  weights[ 4][48]<= -77;  weights[ 4][49]<=  36;  weights[ 4][50]<= 277;  weights[ 4][51]<= 135;  weights[ 4][52]<= 158;  weights[ 4][53]<=  94;  weights[ 4][54]<=-304;  weights[ 4][55]<= 164;  weights[ 4][56]<=  22;  weights[ 4][57]<=  17;  weights[ 4][58]<=  32;  weights[ 4][59]<=-177;  
        weights[ 5][0]<=-200;  weights[ 5][1]<= 106;  weights[ 5][2]<= 288;  weights[ 5][3]<= -96;  weights[ 5][4]<=-155;  weights[ 5][5]<= -46;  weights[ 5][6]<=  22;  weights[ 5][7]<=-239;  weights[ 5][8]<=-214;  weights[ 5][9]<= -10;  weights[ 5][10]<=-265;  weights[ 5][11]<= -61;  weights[ 5][12]<=-117;  weights[ 5][13]<= -34;  weights[ 5][14]<=-127;  weights[ 5][15]<=  22;  weights[ 5][16]<=-159;  weights[ 5][17]<=  51;  weights[ 5][18]<=   7;  weights[ 5][19]<=   6;  weights[ 5][20]<= -36;  weights[ 5][21]<= 245;  weights[ 5][22]<=  62;  weights[ 5][23]<=-142;  weights[ 5][24]<=-130;  weights[ 5][25]<= -41;  weights[ 5][26]<= -10;  weights[ 5][27]<= -12;  weights[ 5][28]<=-107;  weights[ 5][29]<= -65;  weights[ 5][30]<=-113;  weights[ 5][31]<=-175;  weights[ 5][32]<=-123;  weights[ 5][33]<= 248;  weights[ 5][34]<= 108;  weights[ 5][35]<= 127;  weights[ 5][36]<=-285;  weights[ 5][37]<= 153;  weights[ 5][38]<=   6;  weights[ 5][39]<=  31;  weights[ 5][40]<=  19;  weights[ 5][41]<=-164;  weights[ 5][42]<=-107;  weights[ 5][43]<=  27;  weights[ 5][44]<= -51;  weights[ 5][45]<= -53;  weights[ 5][46]<= 144;  weights[ 5][47]<=  71;  weights[ 5][48]<=-164;  weights[ 5][49]<= -20;  weights[ 5][50]<=  47;  weights[ 5][51]<= 240;  weights[ 5][52]<= 285;  weights[ 5][53]<=-151;  weights[ 5][54]<=-288;  weights[ 5][55]<=  83;  weights[ 5][56]<= -67;  weights[ 5][57]<=  43;  weights[ 5][58]<= 332;  weights[ 5][59]<=-199;  
        weights[ 6][0]<=  98;  weights[ 6][1]<= -85;  weights[ 6][2]<=  15;  weights[ 6][3]<=-280;  weights[ 6][4]<= 154;  weights[ 6][5]<= 126;  weights[ 6][6]<=-178;  weights[ 6][7]<= -70;  weights[ 6][8]<=   3;  weights[ 6][9]<=-106;  weights[ 6][10]<=-195;  weights[ 6][11]<=-124;  weights[ 6][12]<=-214;  weights[ 6][13]<=-135;  weights[ 6][14]<=-154;  weights[ 6][15]<=  26;  weights[ 6][16]<= 109;  weights[ 6][17]<=-139;  weights[ 6][18]<=   3;  weights[ 6][19]<=  50;  weights[ 6][20]<=  32;  weights[ 6][21]<= -16;  weights[ 6][22]<=-136;  weights[ 6][23]<= 108;  weights[ 6][24]<=  29;  weights[ 6][25]<=-266;  weights[ 6][26]<= 253;  weights[ 6][27]<=  81;  weights[ 6][28]<=-229;  weights[ 6][29]<= -98;  weights[ 6][30]<= -85;  weights[ 6][31]<= -72;  weights[ 6][32]<= -95;  weights[ 6][33]<= -53;  weights[ 6][34]<=-120;  weights[ 6][35]<=-252;  weights[ 6][36]<= 155;  weights[ 6][37]<= 184;  weights[ 6][38]<=-105;  weights[ 6][39]<=  94;  weights[ 6][40]<= -90;  weights[ 6][41]<=  52;  weights[ 6][42]<= 123;  weights[ 6][43]<=-256;  weights[ 6][44]<=-295;  weights[ 6][45]<=-238;  weights[ 6][46]<= 195;  weights[ 6][47]<= -33;  weights[ 6][48]<= 251;  weights[ 6][49]<=  62;  weights[ 6][50]<=  11;  weights[ 6][51]<= 107;  weights[ 6][52]<= 175;  weights[ 6][53]<=-117;  weights[ 6][54]<= 124;  weights[ 6][55]<=  -3;  weights[ 6][56]<= -74;  weights[ 6][57]<= 221;  weights[ 6][58]<=  29;  weights[ 6][59]<=  43;  
        weights[ 7][0]<= 257;  weights[ 7][1]<=-117;  weights[ 7][2]<=   0;  weights[ 7][3]<=-203;  weights[ 7][4]<= -50;  weights[ 7][5]<= 200;  weights[ 7][6]<=-185;  weights[ 7][7]<=  -1;  weights[ 7][8]<= 171;  weights[ 7][9]<=-141;  weights[ 7][10]<= -16;  weights[ 7][11]<=   3;  weights[ 7][12]<= -62;  weights[ 7][13]<=-111;  weights[ 7][14]<=-163;  weights[ 7][15]<=  -6;  weights[ 7][16]<=-161;  weights[ 7][17]<= 137;  weights[ 7][18]<=-214;  weights[ 7][19]<= -66;  weights[ 7][20]<= -12;  weights[ 7][21]<= 256;  weights[ 7][22]<=  23;  weights[ 7][23]<=  91;  weights[ 7][24]<=-196;  weights[ 7][25]<= -16;  weights[ 7][26]<=-184;  weights[ 7][27]<= 134;  weights[ 7][28]<= -97;  weights[ 7][29]<= 183;  weights[ 7][30]<= 245;  weights[ 7][31]<= 157;  weights[ 7][32]<=-139;  weights[ 7][33]<=-333;  weights[ 7][34]<= -81;  weights[ 7][35]<= -41;  weights[ 7][36]<= 123;  weights[ 7][37]<=-130;  weights[ 7][38]<= 161;  weights[ 7][39]<=-125;  weights[ 7][40]<= 142;  weights[ 7][41]<= 102;  weights[ 7][42]<=-118;  weights[ 7][43]<= -39;  weights[ 7][44]<=-255;  weights[ 7][45]<=  80;  weights[ 7][46]<=  70;  weights[ 7][47]<= 187;  weights[ 7][48]<=-154;  weights[ 7][49]<= -21;  weights[ 7][50]<= 228;  weights[ 7][51]<= -44;  weights[ 7][52]<=-115;  weights[ 7][53]<=  97;  weights[ 7][54]<= -61;  weights[ 7][55]<=-134;  weights[ 7][56]<=  40;  weights[ 7][57]<= 234;  weights[ 7][58]<= 169;  weights[ 7][59]<=-158;  
        weights[ 8][0]<= -14;  weights[ 8][1]<=-268;  weights[ 8][2]<=  23;  weights[ 8][3]<=-209;  weights[ 8][4]<= 200;  weights[ 8][5]<=  80;  weights[ 8][6]<=-176;  weights[ 8][7]<=  49;  weights[ 8][8]<= 115;  weights[ 8][9]<=-113;  weights[ 8][10]<= 204;  weights[ 8][11]<=-156;  weights[ 8][12]<= 108;  weights[ 8][13]<=  78;  weights[ 8][14]<=-113;  weights[ 8][15]<=-215;  weights[ 8][16]<=  74;  weights[ 8][17]<= 199;  weights[ 8][18]<= -67;  weights[ 8][19]<=  97;  weights[ 8][20]<=-138;  weights[ 8][21]<= 241;  weights[ 8][22]<=  85;  weights[ 8][23]<=-147;  weights[ 8][24]<= -55;  weights[ 8][25]<=-159;  weights[ 8][26]<=  99;  weights[ 8][27]<=-216;  weights[ 8][28]<=-159;  weights[ 8][29]<=  42;  weights[ 8][30]<= 103;  weights[ 8][31]<= 207;  weights[ 8][32]<= 200;  weights[ 8][33]<=  75;  weights[ 8][34]<= -42;  weights[ 8][35]<=-210;  weights[ 8][36]<= 137;  weights[ 8][37]<=-121;  weights[ 8][38]<= -20;  weights[ 8][39]<= 107;  weights[ 8][40]<= 204;  weights[ 8][41]<= -95;  weights[ 8][42]<=-208;  weights[ 8][43]<=-101;  weights[ 8][44]<=  50;  weights[ 8][45]<=-175;  weights[ 8][46]<=  53;  weights[ 8][47]<=-126;  weights[ 8][48]<= -79;  weights[ 8][49]<=-206;  weights[ 8][50]<= 252;  weights[ 8][51]<= 253;  weights[ 8][52]<=  24;  weights[ 8][53]<= -50;  weights[ 8][54]<= 247;  weights[ 8][55]<=-197;  weights[ 8][56]<= -89;  weights[ 8][57]<=-171;  weights[ 8][58]<= 187;  weights[ 8][59]<= 293;  
        weights[ 9][0]<= 206;  weights[ 9][1]<=   7;  weights[ 9][2]<=  26;  weights[ 9][3]<=  96;  weights[ 9][4]<= -41;  weights[ 9][5]<=-169;  weights[ 9][6]<=-170;  weights[ 9][7]<= -35;  weights[ 9][8]<= 137;  weights[ 9][9]<= 120;  weights[ 9][10]<=-188;  weights[ 9][11]<=   5;  weights[ 9][12]<= -50;  weights[ 9][13]<= 133;  weights[ 9][14]<=  41;  weights[ 9][15]<=-181;  weights[ 9][16]<=-231;  weights[ 9][17]<= 250;  weights[ 9][18]<=-252;  weights[ 9][19]<= -24;  weights[ 9][20]<=-266;  weights[ 9][21]<= -81;  weights[ 9][22]<=-187;  weights[ 9][23]<= -86;  weights[ 9][24]<=-169;  weights[ 9][25]<= -84;  weights[ 9][26]<= 244;  weights[ 9][27]<=  -1;  weights[ 9][28]<=  40;  weights[ 9][29]<=  38;  weights[ 9][30]<= 190;  weights[ 9][31]<= 229;  weights[ 9][32]<=  71;  weights[ 9][33]<= 148;  weights[ 9][34]<= -48;  weights[ 9][35]<= -21;  weights[ 9][36]<= 209;  weights[ 9][37]<= -48;  weights[ 9][38]<=  -7;  weights[ 9][39]<= 174;  weights[ 9][40]<= -87;  weights[ 9][41]<=-310;  weights[ 9][42]<=  91;  weights[ 9][43]<= -84;  weights[ 9][44]<= 197;  weights[ 9][45]<=  22;  weights[ 9][46]<= 235;  weights[ 9][47]<=  -8;  weights[ 9][48]<= -79;  weights[ 9][49]<=  80;  weights[ 9][50]<= 178;  weights[ 9][51]<=-183;  weights[ 9][52]<= 201;  weights[ 9][53]<= -63;  weights[ 9][54]<=-117;  weights[ 9][55]<=-134;  weights[ 9][56]<= -41;  weights[ 9][57]<=  46;  weights[ 9][58]<= -63;  weights[ 9][59]<= 193;  
        weights[10][0]<=-180;  weights[10][1]<= 178;  weights[10][2]<= -76;  weights[10][3]<=-105;  weights[10][4]<=-197;  weights[10][5]<= 179;  weights[10][6]<=-116;  weights[10][7]<= -31;  weights[10][8]<=-212;  weights[10][9]<=  61;  weights[10][10]<= -96;  weights[10][11]<=-207;  weights[10][12]<= 107;  weights[10][13]<=-277;  weights[10][14]<=-186;  weights[10][15]<= 168;  weights[10][16]<=   5;  weights[10][17]<= 175;  weights[10][18]<= -31;  weights[10][19]<= 164;  weights[10][20]<= 250;  weights[10][21]<=-131;  weights[10][22]<= 132;  weights[10][23]<=  67;  weights[10][24]<=  47;  weights[10][25]<= -46;  weights[10][26]<=  30;  weights[10][27]<= 233;  weights[10][28]<= -25;  weights[10][29]<= -26;  weights[10][30]<=-180;  weights[10][31]<= 205;  weights[10][32]<=  27;  weights[10][33]<= -17;  weights[10][34]<=-177;  weights[10][35]<= 288;  weights[10][36]<=  -4;  weights[10][37]<= 146;  weights[10][38]<=-101;  weights[10][39]<=-169;  weights[10][40]<=  59;  weights[10][41]<=  50;  weights[10][42]<=-164;  weights[10][43]<=-174;  weights[10][44]<=-195;  weights[10][45]<= 242;  weights[10][46]<= 225;  weights[10][47]<= -73;  weights[10][48]<=-231;  weights[10][49]<= -74;  weights[10][50]<=-123;  weights[10][51]<= 243;  weights[10][52]<= -84;  weights[10][53]<=  79;  weights[10][54]<= 246;  weights[10][55]<=-181;  weights[10][56]<= -68;  weights[10][57]<= -11;  weights[10][58]<= 123;  weights[10][59]<= 248;  
        weights[11][0]<= 113;  weights[11][1]<=  33;  weights[11][2]<= -44;  weights[11][3]<= -69;  weights[11][4]<=  92;  weights[11][5]<=-155;  weights[11][6]<= 204;  weights[11][7]<=-110;  weights[11][8]<=-276;  weights[11][9]<=-219;  weights[11][10]<= 170;  weights[11][11]<= 154;  weights[11][12]<=-196;  weights[11][13]<=  71;  weights[11][14]<=-166;  weights[11][15]<=-146;  weights[11][16]<= -58;  weights[11][17]<= 268;  weights[11][18]<=  -4;  weights[11][19]<=  60;  weights[11][20]<=  81;  weights[11][21]<=-187;  weights[11][22]<= -51;  weights[11][23]<=  23;  weights[11][24]<= 142;  weights[11][25]<=-170;  weights[11][26]<= -14;  weights[11][27]<=-179;  weights[11][28]<=  62;  weights[11][29]<=-139;  weights[11][30]<= 173;  weights[11][31]<=-208;  weights[11][32]<= 183;  weights[11][33]<= -28;  weights[11][34]<= -10;  weights[11][35]<= 191;  weights[11][36]<=  51;  weights[11][37]<= -64;  weights[11][38]<=  87;  weights[11][39]<= 110;  weights[11][40]<= 237;  weights[11][41]<=  47;  weights[11][42]<= 247;  weights[11][43]<=-171;  weights[11][44]<=-168;  weights[11][45]<= 116;  weights[11][46]<= -23;  weights[11][47]<=   0;  weights[11][48]<= -99;  weights[11][49]<= -53;  weights[11][50]<= 154;  weights[11][51]<=-108;  weights[11][52]<=  37;  weights[11][53]<=-227;  weights[11][54]<=-111;  weights[11][55]<= -56;  weights[11][56]<=-214;  weights[11][57]<= -78;  weights[11][58]<=  38;  weights[11][59]<= -67;  
        weights[12][0]<= 195;  weights[12][1]<=-171;  weights[12][2]<= 220;  weights[12][3]<=  82;  weights[12][4]<= 205;  weights[12][5]<= 173;  weights[12][6]<= 156;  weights[12][7]<=-243;  weights[12][8]<=-185;  weights[12][9]<= -38;  weights[12][10]<= -84;  weights[12][11]<= 191;  weights[12][12]<=-197;  weights[12][13]<=  63;  weights[12][14]<=-196;  weights[12][15]<=-297;  weights[12][16]<=-210;  weights[12][17]<= -88;  weights[12][18]<=-118;  weights[12][19]<= -54;  weights[12][20]<= 131;  weights[12][21]<= 248;  weights[12][22]<=-128;  weights[12][23]<=-144;  weights[12][24]<=   6;  weights[12][25]<=-134;  weights[12][26]<= 239;  weights[12][27]<=-122;  weights[12][28]<= 123;  weights[12][29]<=  37;  weights[12][30]<=-275;  weights[12][31]<= 165;  weights[12][32]<= 145;  weights[12][33]<=-120;  weights[12][34]<=  54;  weights[12][35]<= 151;  weights[12][36]<= -48;  weights[12][37]<= 227;  weights[12][38]<=  55;  weights[12][39]<= -54;  weights[12][40]<=-167;  weights[12][41]<= 183;  weights[12][42]<=  59;  weights[12][43]<= -48;  weights[12][44]<=-366;  weights[12][45]<=  50;  weights[12][46]<=-239;  weights[12][47]<=  18;  weights[12][48]<= -15;  weights[12][49]<= 155;  weights[12][50]<=-264;  weights[12][51]<=-447;  weights[12][52]<= 193;  weights[12][53]<=-120;  weights[12][54]<=-207;  weights[12][55]<= 241;  weights[12][56]<=-139;  weights[12][57]<= 149;  weights[12][58]<= -72;  weights[12][59]<=-247;  
        weights[13][0]<=-186;  weights[13][1]<=  77;  weights[13][2]<= -38;  weights[13][3]<= -14;  weights[13][4]<= -33;  weights[13][5]<=-143;  weights[13][6]<= -69;  weights[13][7]<=-148;  weights[13][8]<=-223;  weights[13][9]<= 234;  weights[13][10]<= 176;  weights[13][11]<= 110;  weights[13][12]<=  37;  weights[13][13]<= -87;  weights[13][14]<= -11;  weights[13][15]<=  23;  weights[13][16]<=  60;  weights[13][17]<=-115;  weights[13][18]<= -40;  weights[13][19]<= -90;  weights[13][20]<= -49;  weights[13][21]<= -37;  weights[13][22]<=  64;  weights[13][23]<=-145;  weights[13][24]<=-169;  weights[13][25]<= 172;  weights[13][26]<= -13;  weights[13][27]<= 118;  weights[13][28]<= -26;  weights[13][29]<=-121;  weights[13][30]<=  64;  weights[13][31]<=-188;  weights[13][32]<=-204;  weights[13][33]<= 159;  weights[13][34]<= 117;  weights[13][35]<=  56;  weights[13][36]<=-197;  weights[13][37]<= 128;  weights[13][38]<= -19;  weights[13][39]<=-105;  weights[13][40]<=-120;  weights[13][41]<=-135;  weights[13][42]<=-132;  weights[13][43]<= 141;  weights[13][44]<= 141;  weights[13][45]<= -78;  weights[13][46]<=-203;  weights[13][47]<= 177;  weights[13][48]<= 201;  weights[13][49]<=-149;  weights[13][50]<=  39;  weights[13][51]<= 253;  weights[13][52]<= -56;  weights[13][53]<=-157;  weights[13][54]<=  23;  weights[13][55]<=-138;  weights[13][56]<=  80;  weights[13][57]<= -24;  weights[13][58]<= -42;  weights[13][59]<=  88;  
        weights[14][0]<= 244;  weights[14][1]<=   3;  weights[14][2]<=  93;  weights[14][3]<= -99;  weights[14][4]<= 209;  weights[14][5]<= -31;  weights[14][6]<= 162;  weights[14][7]<=-150;  weights[14][8]<=-173;  weights[14][9]<=-163;  weights[14][10]<=  84;  weights[14][11]<=-190;  weights[14][12]<=  74;  weights[14][13]<= 272;  weights[14][14]<= 128;  weights[14][15]<=-104;  weights[14][16]<= 160;  weights[14][17]<= -15;  weights[14][18]<=-172;  weights[14][19]<=  64;  weights[14][20]<=  77;  weights[14][21]<=  85;  weights[14][22]<=  40;  weights[14][23]<= 128;  weights[14][24]<= 264;  weights[14][25]<= -67;  weights[14][26]<= 124;  weights[14][27]<=-309;  weights[14][28]<= -38;  weights[14][29]<= -70;  weights[14][30]<= 207;  weights[14][31]<=-167;  weights[14][32]<= 131;  weights[14][33]<=  45;  weights[14][34]<=  84;  weights[14][35]<= -29;  weights[14][36]<= -89;  weights[14][37]<=  23;  weights[14][38]<=   0;  weights[14][39]<=-187;  weights[14][40]<=-212;  weights[14][41]<=  29;  weights[14][42]<= -47;  weights[14][43]<=-150;  weights[14][44]<=-106;  weights[14][45]<=  70;  weights[14][46]<=-161;  weights[14][47]<= 106;  weights[14][48]<=-168;  weights[14][49]<=  10;  weights[14][50]<=  46;  weights[14][51]<=-116;  weights[14][52]<= 160;  weights[14][53]<= -46;  weights[14][54]<= 181;  weights[14][55]<=-194;  weights[14][56]<=  69;  weights[14][57]<=  23;  weights[14][58]<=-182;  weights[14][59]<= 136;  
        weights[15][0]<=-235;  weights[15][1]<=  56;  weights[15][2]<=  38;  weights[15][3]<=  20;  weights[15][4]<=-256;  weights[15][5]<= -58;  weights[15][6]<=-239;  weights[15][7]<= 152;  weights[15][8]<=  79;  weights[15][9]<=  95;  weights[15][10]<= -46;  weights[15][11]<= -64;  weights[15][12]<= -78;  weights[15][13]<=  46;  weights[15][14]<=-140;  weights[15][15]<=-150;  weights[15][16]<=-217;  weights[15][17]<=   2;  weights[15][18]<=-225;  weights[15][19]<=  19;  weights[15][20]<=  38;  weights[15][21]<= 178;  weights[15][22]<= -55;  weights[15][23]<= 116;  weights[15][24]<=  59;  weights[15][25]<= -78;  weights[15][26]<= 100;  weights[15][27]<= 129;  weights[15][28]<= -98;  weights[15][29]<=  26;  weights[15][30]<=-160;  weights[15][31]<=  -9;  weights[15][32]<= 140;  weights[15][33]<= -26;  weights[15][34]<=  -1;  weights[15][35]<=-142;  weights[15][36]<= -13;  weights[15][37]<=   8;  weights[15][38]<=-144;  weights[15][39]<= 114;  weights[15][40]<=-139;  weights[15][41]<=-113;  weights[15][42]<= 232;  weights[15][43]<=  42;  weights[15][44]<= 146;  weights[15][45]<=-258;  weights[15][46]<=-173;  weights[15][47]<= 232;  weights[15][48]<= -13;  weights[15][49]<=-147;  weights[15][50]<=-199;  weights[15][51]<= 191;  weights[15][52]<=-126;  weights[15][53]<=  20;  weights[15][54]<=  99;  weights[15][55]<=  33;  weights[15][56]<=-193;  weights[15][57]<= 193;  weights[15][58]<= 264;  weights[15][59]<= 194;  
        weights[16][0]<= 257;  weights[16][1]<=-206;  weights[16][2]<=-201;  weights[16][3]<= 219;  weights[16][4]<=-112;  weights[16][5]<= -34;  weights[16][6]<= -60;  weights[16][7]<=-137;  weights[16][8]<=-132;  weights[16][9]<=  -1;  weights[16][10]<=  88;  weights[16][11]<= 189;  weights[16][12]<= -59;  weights[16][13]<= -33;  weights[16][14]<= -86;  weights[16][15]<=  87;  weights[16][16]<=-244;  weights[16][17]<= 226;  weights[16][18]<= 267;  weights[16][19]<=  20;  weights[16][20]<= 279;  weights[16][21]<= -38;  weights[16][22]<= 259;  weights[16][23]<=-111;  weights[16][24]<=  -1;  weights[16][25]<= 122;  weights[16][26]<=  74;  weights[16][27]<=-272;  weights[16][28]<= 191;  weights[16][29]<= 128;  weights[16][30]<= 214;  weights[16][31]<=-169;  weights[16][32]<=-139;  weights[16][33]<= 103;  weights[16][34]<= -65;  weights[16][35]<=-137;  weights[16][36]<=-194;  weights[16][37]<=-171;  weights[16][38]<= -70;  weights[16][39]<=-220;  weights[16][40]<= -50;  weights[16][41]<=  76;  weights[16][42]<=-176;  weights[16][43]<= 138;  weights[16][44]<= -11;  weights[16][45]<=  88;  weights[16][46]<=   0;  weights[16][47]<= 120;  weights[16][48]<=-189;  weights[16][49]<= -93;  weights[16][50]<= 163;  weights[16][51]<= 243;  weights[16][52]<=  82;  weights[16][53]<=  98;  weights[16][54]<= 149;  weights[16][55]<=-199;  weights[16][56]<=-136;  weights[16][57]<= -46;  weights[16][58]<=-184;  weights[16][59]<= 223;  
        weights[17][0]<=-206;  weights[17][1]<=-197;  weights[17][2]<=-294;  weights[17][3]<= 141;  weights[17][4]<=  12;  weights[17][5]<= 115;  weights[17][6]<= 237;  weights[17][7]<=  74;  weights[17][8]<= -44;  weights[17][9]<=-131;  weights[17][10]<= 228;  weights[17][11]<= 196;  weights[17][12]<= 172;  weights[17][13]<=  14;  weights[17][14]<=  77;  weights[17][15]<=  29;  weights[17][16]<= -62;  weights[17][17]<= 200;  weights[17][18]<= -38;  weights[17][19]<= -23;  weights[17][20]<= 133;  weights[17][21]<=  -3;  weights[17][22]<= 128;  weights[17][23]<= -97;  weights[17][24]<= 173;  weights[17][25]<= 104;  weights[17][26]<= -91;  weights[17][27]<= -10;  weights[17][28]<= 187;  weights[17][29]<= -76;  weights[17][30]<= -91;  weights[17][31]<=  46;  weights[17][32]<= -33;  weights[17][33]<=-242;  weights[17][34]<= -32;  weights[17][35]<= 181;  weights[17][36]<=  85;  weights[17][37]<=-186;  weights[17][38]<= -98;  weights[17][39]<= -53;  weights[17][40]<=-191;  weights[17][41]<=  31;  weights[17][42]<= -24;  weights[17][43]<=  63;  weights[17][44]<= -11;  weights[17][45]<=-189;  weights[17][46]<=-232;  weights[17][47]<= -40;  weights[17][48]<=  70;  weights[17][49]<= 140;  weights[17][50]<= -16;  weights[17][51]<=-279;  weights[17][52]<=  73;  weights[17][53]<= 158;  weights[17][54]<= 105;  weights[17][55]<= 181;  weights[17][56]<=  46;  weights[17][57]<= -22;  weights[17][58]<=  18;  weights[17][59]<=-105;  
        weights[18][0]<= 131;  weights[18][1]<=-208;  weights[18][2]<= 139;  weights[18][3]<=-188;  weights[18][4]<=-101;  weights[18][5]<= -22;  weights[18][6]<=  80;  weights[18][7]<= 121;  weights[18][8]<=-235;  weights[18][9]<= -99;  weights[18][10]<= -15;  weights[18][11]<=  78;  weights[18][12]<=  87;  weights[18][13]<=-138;  weights[18][14]<=  24;  weights[18][15]<=-176;  weights[18][16]<=   2;  weights[18][17]<=  67;  weights[18][18]<=-213;  weights[18][19]<= -81;  weights[18][20]<= 111;  weights[18][21]<=  38;  weights[18][22]<=-239;  weights[18][23]<=  62;  weights[18][24]<= -12;  weights[18][25]<= 126;  weights[18][26]<= -24;  weights[18][27]<= 117;  weights[18][28]<= 118;  weights[18][29]<= 108;  weights[18][30]<= 132;  weights[18][31]<= 153;  weights[18][32]<= 151;  weights[18][33]<= 159;  weights[18][34]<= 142;  weights[18][35]<= 227;  weights[18][36]<=-153;  weights[18][37]<= -16;  weights[18][38]<= -77;  weights[18][39]<=  14;  weights[18][40]<= 113;  weights[18][41]<= -44;  weights[18][42]<=  68;  weights[18][43]<= -71;  weights[18][44]<=-289;  weights[18][45]<= 142;  weights[18][46]<= -88;  weights[18][47]<=  11;  weights[18][48]<= 180;  weights[18][49]<= -55;  weights[18][50]<=-183;  weights[18][51]<=  20;  weights[18][52]<=  92;  weights[18][53]<= 155;  weights[18][54]<=  41;  weights[18][55]<= 162;  weights[18][56]<=-186;  weights[18][57]<=-194;  weights[18][58]<= 167;  weights[18][59]<=-115;  
        weights[19][0]<= -19;  weights[19][1]<= 111;  weights[19][2]<=  11;  weights[19][3]<= -95;  weights[19][4]<=-196;  weights[19][5]<=-125;  weights[19][6]<= 278;  weights[19][7]<=  97;  weights[19][8]<=  25;  weights[19][9]<=  20;  weights[19][10]<=-140;  weights[19][11]<= -78;  weights[19][12]<= 124;  weights[19][13]<=-200;  weights[19][14]<=  25;  weights[19][15]<= 120;  weights[19][16]<=-158;  weights[19][17]<=-120;  weights[19][18]<= -70;  weights[19][19]<= -16;  weights[19][20]<=  99;  weights[19][21]<=-142;  weights[19][22]<=  66;  weights[19][23]<=-178;  weights[19][24]<=  88;  weights[19][25]<=  52;  weights[19][26]<= 108;  weights[19][27]<=  -4;  weights[19][28]<=  91;  weights[19][29]<=-117;  weights[19][30]<=-179;  weights[19][31]<= 149;  weights[19][32]<=-132;  weights[19][33]<=  -3;  weights[19][34]<= -96;  weights[19][35]<=  73;  weights[19][36]<=-227;  weights[19][37]<=  51;  weights[19][38]<= 112;  weights[19][39]<= 144;  weights[19][40]<=  69;  weights[19][41]<= 110;  weights[19][42]<= 206;  weights[19][43]<=-201;  weights[19][44]<=-325;  weights[19][45]<= 245;  weights[19][46]<= -65;  weights[19][47]<=  60;  weights[19][48]<= 109;  weights[19][49]<= 221;  weights[19][50]<= -41;  weights[19][51]<=-114;  weights[19][52]<= 131;  weights[19][53]<=  50;  weights[19][54]<= 245;  weights[19][55]<=-131;  weights[19][56]<= 130;  weights[19][57]<= 199;  weights[19][58]<= 142;  weights[19][59]<=-351;  
        weights[20][0]<=-110;  weights[20][1]<= 173;  weights[20][2]<=-114;  weights[20][3]<= 170;  weights[20][4]<=  44;  weights[20][5]<= -51;  weights[20][6]<=-167;  weights[20][7]<= -89;  weights[20][8]<=-186;  weights[20][9]<=  64;  weights[20][10]<= 234;  weights[20][11]<=-281;  weights[20][12]<= 152;  weights[20][13]<= -95;  weights[20][14]<= 231;  weights[20][15]<=  -1;  weights[20][16]<=  56;  weights[20][17]<= 129;  weights[20][18]<= -42;  weights[20][19]<= -88;  weights[20][20]<= 249;  weights[20][21]<= -19;  weights[20][22]<=  62;  weights[20][23]<= -28;  weights[20][24]<= 223;  weights[20][25]<=-274;  weights[20][26]<= 128;  weights[20][27]<=-169;  weights[20][28]<=  18;  weights[20][29]<=  40;  weights[20][30]<=  17;  weights[20][31]<=-188;  weights[20][32]<=  99;  weights[20][33]<=  68;  weights[20][34]<= -20;  weights[20][35]<= 157;  weights[20][36]<=-142;  weights[20][37]<= 116;  weights[20][38]<=  82;  weights[20][39]<=-290;  weights[20][40]<=-139;  weights[20][41]<=-118;  weights[20][42]<=  49;  weights[20][43]<=  52;  weights[20][44]<=  80;  weights[20][45]<= 195;  weights[20][46]<=-216;  weights[20][47]<=-171;  weights[20][48]<=-192;  weights[20][49]<=-139;  weights[20][50]<=  30;  weights[20][51]<= 267;  weights[20][52]<=-143;  weights[20][53]<= 165;  weights[20][54]<= 127;  weights[20][55]<=-133;  weights[20][56]<=  19;  weights[20][57]<=-197;  weights[20][58]<= -56;  weights[20][59]<=  94;  
        weights[21][0]<=-171;  weights[21][1]<= -78;  weights[21][2]<=  97;  weights[21][3]<= -30;  weights[21][4]<=-116;  weights[21][5]<=  14;  weights[21][6]<=-198;  weights[21][7]<= -85;  weights[21][8]<= 257;  weights[21][9]<= 158;  weights[21][10]<=-186;  weights[21][11]<= -36;  weights[21][12]<= 234;  weights[21][13]<= -79;  weights[21][14]<= 202;  weights[21][15]<=-150;  weights[21][16]<=  70;  weights[21][17]<= -85;  weights[21][18]<= 137;  weights[21][19]<=  71;  weights[21][20]<=-142;  weights[21][21]<= -82;  weights[21][22]<= 128;  weights[21][23]<=  32;  weights[21][24]<=-110;  weights[21][25]<= 103;  weights[21][26]<=-117;  weights[21][27]<= 201;  weights[21][28]<=-235;  weights[21][29]<= -49;  weights[21][30]<= 123;  weights[21][31]<=  75;  weights[21][32]<=-155;  weights[21][33]<= 242;  weights[21][34]<= -59;  weights[21][35]<= 130;  weights[21][36]<= 218;  weights[21][37]<= -35;  weights[21][38]<= -99;  weights[21][39]<=  69;  weights[21][40]<=-170;  weights[21][41]<= -29;  weights[21][42]<= -48;  weights[21][43]<= -21;  weights[21][44]<= 173;  weights[21][45]<=   1;  weights[21][46]<=-105;  weights[21][47]<=-110;  weights[21][48]<= 213;  weights[21][49]<= 120;  weights[21][50]<= 193;  weights[21][51]<=-225;  weights[21][52]<=  36;  weights[21][53]<= 119;  weights[21][54]<=  61;  weights[21][55]<= -11;  weights[21][56]<=-186;  weights[21][57]<= -68;  weights[21][58]<=-109;  weights[21][59]<=-172;  
        weights[22][0]<=-117;  weights[22][1]<=  70;  weights[22][2]<= -43;  weights[22][3]<= 304;  weights[22][4]<=-103;  weights[22][5]<= 239;  weights[22][6]<=-164;  weights[22][7]<= 109;  weights[22][8]<=-197;  weights[22][9]<=-176;  weights[22][10]<=-138;  weights[22][11]<=  23;  weights[22][12]<= -97;  weights[22][13]<= -81;  weights[22][14]<=  64;  weights[22][15]<=-210;  weights[22][16]<=  51;  weights[22][17]<= 220;  weights[22][18]<=-145;  weights[22][19]<=-221;  weights[22][20]<=-285;  weights[22][21]<= 101;  weights[22][22]<=  18;  weights[22][23]<=  26;  weights[22][24]<=  90;  weights[22][25]<= 279;  weights[22][26]<=-119;  weights[22][27]<= -40;  weights[22][28]<=-167;  weights[22][29]<= 119;  weights[22][30]<= 138;  weights[22][31]<=  95;  weights[22][32]<=   1;  weights[22][33]<= 295;  weights[22][34]<= 187;  weights[22][35]<= -65;  weights[22][36]<= 332;  weights[22][37]<= -65;  weights[22][38]<= -35;  weights[22][39]<= 111;  weights[22][40]<=-176;  weights[22][41]<= 234;  weights[22][42]<= -35;  weights[22][43]<=  56;  weights[22][44]<= 233;  weights[22][45]<=-209;  weights[22][46]<= 111;  weights[22][47]<= -49;  weights[22][48]<=-107;  weights[22][49]<= 127;  weights[22][50]<=-187;  weights[22][51]<= 128;  weights[22][52]<=   3;  weights[22][53]<= -97;  weights[22][54]<=  80;  weights[22][55]<=-212;  weights[22][56]<= -48;  weights[22][57]<= -78;  weights[22][58]<= -95;  weights[22][59]<= 209;  
        weights[23][0]<= 121;  weights[23][1]<=  42;  weights[23][2]<= 214;  weights[23][3]<=-100;  weights[23][4]<=-119;  weights[23][5]<= 105;  weights[23][6]<= -97;  weights[23][7]<=-121;  weights[23][8]<= 176;  weights[23][9]<= 293;  weights[23][10]<=-116;  weights[23][11]<= 105;  weights[23][12]<= -92;  weights[23][13]<=-137;  weights[23][14]<=-194;  weights[23][15]<=-117;  weights[23][16]<= 247;  weights[23][17]<=-199;  weights[23][18]<= 127;  weights[23][19]<=  70;  weights[23][20]<=-165;  weights[23][21]<= -27;  weights[23][22]<= -88;  weights[23][23]<=-120;  weights[23][24]<=-191;  weights[23][25]<= -45;  weights[23][26]<= -35;  weights[23][27]<=-115;  weights[23][28]<=  13;  weights[23][29]<= 114;  weights[23][30]<=-181;  weights[23][31]<= 103;  weights[23][32]<=-169;  weights[23][33]<=  64;  weights[23][34]<=   2;  weights[23][35]<=  70;  weights[23][36]<=-140;  weights[23][37]<=  23;  weights[23][38]<= 201;  weights[23][39]<= 172;  weights[23][40]<= -33;  weights[23][41]<=-252;  weights[23][42]<=-122;  weights[23][43]<=-116;  weights[23][44]<= -11;  weights[23][45]<=  54;  weights[23][46]<= 247;  weights[23][47]<= 164;  weights[23][48]<= 247;  weights[23][49]<=-114;  weights[23][50]<=-222;  weights[23][51]<= 210;  weights[23][52]<= 250;  weights[23][53]<=-211;  weights[23][54]<= -74;  weights[23][55]<= -91;  weights[23][56]<=   8;  weights[23][57]<= 167;  weights[23][58]<= -71;  weights[23][59]<= 194;  
        weights[24][0]<= 164;  weights[24][1]<=-179;  weights[24][2]<=-175;  weights[24][3]<=  34;  weights[24][4]<=-135;  weights[24][5]<=-150;  weights[24][6]<= -94;  weights[24][7]<=-207;  weights[24][8]<= -13;  weights[24][9]<=  58;  weights[24][10]<= -71;  weights[24][11]<=-100;  weights[24][12]<=  16;  weights[24][13]<=-214;  weights[24][14]<=  42;  weights[24][15]<= -22;  weights[24][16]<=-151;  weights[24][17]<=  75;  weights[24][18]<=   5;  weights[24][19]<= -42;  weights[24][20]<=-204;  weights[24][21]<=-197;  weights[24][22]<=-128;  weights[24][23]<= 327;  weights[24][24]<= 158;  weights[24][25]<=   6;  weights[24][26]<= 111;  weights[24][27]<=-183;  weights[24][28]<= 330;  weights[24][29]<= -48;  weights[24][30]<=-111;  weights[24][31]<=-117;  weights[24][32]<=-130;  weights[24][33]<= -42;  weights[24][34]<= 255;  weights[24][35]<= 126;  weights[24][36]<=  36;  weights[24][37]<=  -6;  weights[24][38]<= -57;  weights[24][39]<= -59;  weights[24][40]<=-168;  weights[24][41]<=  28;  weights[24][42]<= 220;  weights[24][43]<=-271;  weights[24][44]<= 125;  weights[24][45]<= 219;  weights[24][46]<= 232;  weights[24][47]<= 241;  weights[24][48]<=   0;  weights[24][49]<=  26;  weights[24][50]<= -97;  weights[24][51]<=-393;  weights[24][52]<= 102;  weights[24][53]<=-137;  weights[24][54]<= -49;  weights[24][55]<= -50;  weights[24][56]<=-105;  weights[24][57]<= 187;  weights[24][58]<= -66;  weights[24][59]<=-370;  
        weights[25][0]<=  19;  weights[25][1]<= -21;  weights[25][2]<= 241;  weights[25][3]<=  99;  weights[25][4]<=-228;  weights[25][5]<= -50;  weights[25][6]<= 161;  weights[25][7]<= 108;  weights[25][8]<= 212;  weights[25][9]<=  17;  weights[25][10]<=-224;  weights[25][11]<=-214;  weights[25][12]<=  77;  weights[25][13]<=  94;  weights[25][14]<=  59;  weights[25][15]<= -12;  weights[25][16]<=-112;  weights[25][17]<= -61;  weights[25][18]<= 227;  weights[25][19]<= -36;  weights[25][20]<= -70;  weights[25][21]<= 156;  weights[25][22]<=-108;  weights[25][23]<= -44;  weights[25][24]<=  63;  weights[25][25]<=-126;  weights[25][26]<= 124;  weights[25][27]<= -28;  weights[25][28]<= -91;  weights[25][29]<=  33;  weights[25][30]<= -88;  weights[25][31]<=-150;  weights[25][32]<=-131;  weights[25][33]<= 139;  weights[25][34]<=  63;  weights[25][35]<= 112;  weights[25][36]<=  58;  weights[25][37]<= -39;  weights[25][38]<=  27;  weights[25][39]<=  12;  weights[25][40]<= -66;  weights[25][41]<=-161;  weights[25][42]<= 316;  weights[25][43]<=-124;  weights[25][44]<=-103;  weights[25][45]<=-255;  weights[25][46]<= -28;  weights[25][47]<= -81;  weights[25][48]<= 160;  weights[25][49]<= -60;  weights[25][50]<=  48;  weights[25][51]<=-177;  weights[25][52]<=  29;  weights[25][53]<= -68;  weights[25][54]<=-149;  weights[25][55]<= 199;  weights[25][56]<= -97;  weights[25][57]<=-144;  weights[25][58]<=-155;  weights[25][59]<= 214;  
        weights[26][0]<=-311;  weights[26][1]<=-256;  weights[26][2]<=   2;  weights[26][3]<= 186;  weights[26][4]<= 121;  weights[26][5]<=  21;  weights[26][6]<= 102;  weights[26][7]<=   9;  weights[26][8]<= -92;  weights[26][9]<=-150;  weights[26][10]<=  12;  weights[26][11]<=  43;  weights[26][12]<=-205;  weights[26][13]<=  -3;  weights[26][14]<=  18;  weights[26][15]<=  76;  weights[26][16]<= 145;  weights[26][17]<=  67;  weights[26][18]<= 122;  weights[26][19]<= 104;  weights[26][20]<= -32;  weights[26][21]<=-124;  weights[26][22]<= 158;  weights[26][23]<=-174;  weights[26][24]<= -83;  weights[26][25]<=-199;  weights[26][26]<=  53;  weights[26][27]<= 211;  weights[26][28]<= 103;  weights[26][29]<= -96;  weights[26][30]<= 217;  weights[26][31]<= -58;  weights[26][32]<=-146;  weights[26][33]<= 100;  weights[26][34]<=  19;  weights[26][35]<= -23;  weights[26][36]<=  96;  weights[26][37]<=-263;  weights[26][38]<= -36;  weights[26][39]<=  22;  weights[26][40]<=-175;  weights[26][41]<= -81;  weights[26][42]<= 136;  weights[26][43]<= -75;  weights[26][44]<=-194;  weights[26][45]<= 165;  weights[26][46]<=  90;  weights[26][47]<=  18;  weights[26][48]<=  36;  weights[26][49]<= 121;  weights[26][50]<=  82;  weights[26][51]<=-227;  weights[26][52]<=  96;  weights[26][53]<= 264;  weights[26][54]<=  59;  weights[26][55]<= -18;  weights[26][56]<= -70;  weights[26][57]<=-166;  weights[26][58]<=  11;  weights[26][59]<=   1;  
        weights[27][0]<= 239;  weights[27][1]<= 150;  weights[27][2]<=  95;  weights[27][3]<= 168;  weights[27][4]<= 181;  weights[27][5]<= 268;  weights[27][6]<=-223;  weights[27][7]<=-150;  weights[27][8]<= 225;  weights[27][9]<=-168;  weights[27][10]<= -92;  weights[27][11]<=-239;  weights[27][12]<= 153;  weights[27][13]<= -82;  weights[27][14]<=  10;  weights[27][15]<=  46;  weights[27][16]<=-189;  weights[27][17]<= 118;  weights[27][18]<=-119;  weights[27][19]<= -71;  weights[27][20]<= 151;  weights[27][21]<= 113;  weights[27][22]<= -25;  weights[27][23]<=-155;  weights[27][24]<=  -8;  weights[27][25]<= -21;  weights[27][26]<=  37;  weights[27][27]<=-217;  weights[27][28]<=-145;  weights[27][29]<= 169;  weights[27][30]<= -12;  weights[27][31]<=-124;  weights[27][32]<= 226;  weights[27][33]<= -42;  weights[27][34]<= 147;  weights[27][35]<=   5;  weights[27][36]<= -19;  weights[27][37]<= 144;  weights[27][38]<= -81;  weights[27][39]<= -34;  weights[27][40]<=-288;  weights[27][41]<= 193;  weights[27][42]<= 154;  weights[27][43]<=  82;  weights[27][44]<= -87;  weights[27][45]<=-214;  weights[27][46]<=-119;  weights[27][47]<= 187;  weights[27][48]<=-151;  weights[27][49]<=  50;  weights[27][50]<=-168;  weights[27][51]<=  73;  weights[27][52]<=  49;  weights[27][53]<= 134;  weights[27][54]<=  24;  weights[27][55]<= 190;  weights[27][56]<=-239;  weights[27][57]<= -60;  weights[27][58]<=  28;  weights[27][59]<= 136;  
        weights[28][0]<=-112;  weights[28][1]<=-142;  weights[28][2]<=-238;  weights[28][3]<=  48;  weights[28][4]<=  88;  weights[28][5]<= -81;  weights[28][6]<= -32;  weights[28][7]<= 123;  weights[28][8]<=-314;  weights[28][9]<=-160;  weights[28][10]<= -25;  weights[28][11]<= -38;  weights[28][12]<=  87;  weights[28][13]<=  89;  weights[28][14]<=-112;  weights[28][15]<= -93;  weights[28][16]<= -38;  weights[28][17]<= 108;  weights[28][18]<=-290;  weights[28][19]<= -70;  weights[28][20]<=  35;  weights[28][21]<=-185;  weights[28][22]<=  87;  weights[28][23]<= 205;  weights[28][24]<= -66;  weights[28][25]<= -35;  weights[28][26]<= -18;  weights[28][27]<= 104;  weights[28][28]<=-162;  weights[28][29]<= -74;  weights[28][30]<=  86;  weights[28][31]<= 162;  weights[28][32]<=  61;  weights[28][33]<=-312;  weights[28][34]<=-134;  weights[28][35]<= 121;  weights[28][36]<= -81;  weights[28][37]<=  30;  weights[28][38]<=  98;  weights[28][39]<= -70;  weights[28][40]<= 144;  weights[28][41]<=-121;  weights[28][42]<=-130;  weights[28][43]<=-185;  weights[28][44]<= 191;  weights[28][45]<= 146;  weights[28][46]<=-105;  weights[28][47]<= 141;  weights[28][48]<= 142;  weights[28][49]<= 137;  weights[28][50]<= 115;  weights[28][51]<=-306;  weights[28][52]<= -85;  weights[28][53]<= 167;  weights[28][54]<=   4;  weights[28][55]<=-151;  weights[28][56]<= 220;  weights[28][57]<= 122;  weights[28][58]<=-102;  weights[28][59]<=-299;  
        weights[29][0]<=-137;  weights[29][1]<= -35;  weights[29][2]<=  73;  weights[29][3]<=  95;  weights[29][4]<= 175;  weights[29][5]<=-141;  weights[29][6]<=  98;  weights[29][7]<= 150;  weights[29][8]<= -80;  weights[29][9]<= -78;  weights[29][10]<=-297;  weights[29][11]<=-181;  weights[29][12]<= -55;  weights[29][13]<=  97;  weights[29][14]<=  71;  weights[29][15]<= -85;  weights[29][16]<=-171;  weights[29][17]<= 240;  weights[29][18]<= 270;  weights[29][19]<=-116;  weights[29][20]<=  47;  weights[29][21]<= -35;  weights[29][22]<= 103;  weights[29][23]<=-197;  weights[29][24]<= 132;  weights[29][25]<=-205;  weights[29][26]<= -51;  weights[29][27]<= -82;  weights[29][28]<=  15;  weights[29][29]<= -31;  weights[29][30]<= 164;  weights[29][31]<= 111;  weights[29][32]<=  74;  weights[29][33]<=  63;  weights[29][34]<= 138;  weights[29][35]<= 190;  weights[29][36]<=  68;  weights[29][37]<=  94;  weights[29][38]<=  89;  weights[29][39]<=-129;  weights[29][40]<= 253;  weights[29][41]<=-168;  weights[29][42]<=-201;  weights[29][43]<= -64;  weights[29][44]<= 133;  weights[29][45]<= -84;  weights[29][46]<=-137;  weights[29][47]<=  94;  weights[29][48]<=-226;  weights[29][49]<=  92;  weights[29][50]<=-171;  weights[29][51]<=-279;  weights[29][52]<= 177;  weights[29][53]<= 162;  weights[29][54]<=  47;  weights[29][55]<=-117;  weights[29][56]<= -72;  weights[29][57]<=-185;  weights[29][58]<= 149;  weights[29][59]<=-127;  
        weights[30][0]<=-125;  weights[30][1]<= 232;  weights[30][2]<=  -2;  weights[30][3]<= -95;  weights[30][4]<=-126;  weights[30][5]<=  45;  weights[30][6]<= 163;  weights[30][7]<= -23;  weights[30][8]<= -72;  weights[30][9]<=  48;  weights[30][10]<=-191;  weights[30][11]<= 135;  weights[30][12]<=-109;  weights[30][13]<=  86;  weights[30][14]<= 153;  weights[30][15]<=-332;  weights[30][16]<=-108;  weights[30][17]<=-157;  weights[30][18]<=-186;  weights[30][19]<=-134;  weights[30][20]<=-181;  weights[30][21]<=-179;  weights[30][22]<= 140;  weights[30][23]<=-107;  weights[30][24]<=  18;  weights[30][25]<=  69;  weights[30][26]<=-156;  weights[30][27]<= 269;  weights[30][28]<=-136;  weights[30][29]<=-150;  weights[30][30]<=  48;  weights[30][31]<= -30;  weights[30][32]<= 139;  weights[30][33]<=-195;  weights[30][34]<=-203;  weights[30][35]<=  87;  weights[30][36]<=  98;  weights[30][37]<=-119;  weights[30][38]<=-142;  weights[30][39]<= -71;  weights[30][40]<=  61;  weights[30][41]<= 110;  weights[30][42]<= 116;  weights[30][43]<=-157;  weights[30][44]<=-149;  weights[30][45]<= -59;  weights[30][46]<= 139;  weights[30][47]<=-102;  weights[30][48]<=-189;  weights[30][49]<=  56;  weights[30][50]<= -27;  weights[30][51]<=  -9;  weights[30][52]<= -25;  weights[30][53]<= -12;  weights[30][54]<=  12;  weights[30][55]<=-113;  weights[30][56]<= 263;  weights[30][57]<= 196;  weights[30][58]<= 203;  weights[30][59]<=-197;  
        weights[31][0]<= -95;  weights[31][1]<=-221;  weights[31][2]<= -28;  weights[31][3]<= 155;  weights[31][4]<= -87;  weights[31][5]<=  32;  weights[31][6]<=-130;  weights[31][7]<= 151;  weights[31][8]<=-191;  weights[31][9]<= -25;  weights[31][10]<=-238;  weights[31][11]<= 171;  weights[31][12]<=   0;  weights[31][13]<= 203;  weights[31][14]<=-183;  weights[31][15]<=-130;  weights[31][16]<= -52;  weights[31][17]<= -88;  weights[31][18]<= 135;  weights[31][19]<= 150;  weights[31][20]<=  94;  weights[31][21]<=  50;  weights[31][22]<= 175;  weights[31][23]<= -61;  weights[31][24]<= -81;  weights[31][25]<=  99;  weights[31][26]<= 162;  weights[31][27]<=  40;  weights[31][28]<=-235;  weights[31][29]<= -73;  weights[31][30]<=-148;  weights[31][31]<=  75;  weights[31][32]<=-220;  weights[31][33]<= 115;  weights[31][34]<= -75;  weights[31][35]<= 135;  weights[31][36]<=-275;  weights[31][37]<= 126;  weights[31][38]<=  71;  weights[31][39]<= -26;  weights[31][40]<= 197;  weights[31][41]<= 218;  weights[31][42]<= -76;  weights[31][43]<= -48;  weights[31][44]<= 142;  weights[31][45]<=  45;  weights[31][46]<= 114;  weights[31][47]<= -17;  weights[31][48]<=  37;  weights[31][49]<=  87;  weights[31][50]<=-172;  weights[31][51]<= 157;  weights[31][52]<=  33;  weights[31][53]<=  13;  weights[31][54]<=  48;  weights[31][55]<=  40;  weights[31][56]<=  31;  weights[31][57]<=  26;  weights[31][58]<= -59;  weights[31][59]<=-119; 

        biases[ 0]<= 13637;  biases[ 1]<= 19819;  biases[ 2]<=-59667;  biases[ 3]<= 36143;  biases[ 4]<=-38093;  biases[ 5]<= 37491;  biases[ 6]<= 61100;  biases[ 7]<= 19283;  biases[ 8]<= 50092;  biases[ 9]<=  6236;  biases[10]<=-31489;  biases[11]<= 43860;  biases[12]<= -7430;  biases[13]<=   -18;  biases[14]<=-22899;  biases[15]<=-13377;  biases[16]<=  3406;  biases[17]<=-12774;  biases[18]<=  2312;  biases[19]<=-27712;  biases[20]<=-71924;  biases[21]<=-61095;  biases[22]<= -5993;  biases[23]<=-27534;  biases[24]<= 25367;  biases[25]<= 39074;  biases[26]<=-15747;  biases[27]<=-27113;  biases[28]<= 67387;  biases[29]<= 54720;  biases[30]<= 20034;  biases[31]<= 23520; 
    end

    always@(posedge clk) begin
        if(rst||~start) begin
            w<=0;
            b<=0;
            ready<=0;
        end else if(start) begin
            if(input_pixel_addr<60&&output_pixel_addr<32) begin
                w<=weights[output_pixel_addr][input_pixel_addr];
                if(input_pixel_addr==59) begin
                    b<=biases[output_pixel_addr];
                end else begin
                    b<=0;
                end
                ready<=1;
            end else begin
                w<=0;
                b<=0;
                ready<=0;
            end
        end
    end
endmodule